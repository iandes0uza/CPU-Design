library verilog;
use verilog.vl_types.all;
entity control_unit is
    generic(
        r_s             : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        T0              : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        T1              : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        T2              : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        T3              : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        load_T0         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        load_T1         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        load_T2         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        load_T3         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0);
        load_T4         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1);
        loadi_T0        : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        loadi_T1        : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        loadi_T2        : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        store_T0        : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        store_T1        : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1);
        store_T2        : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        store_T3        : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1);
        alu2_T0         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0);
        alu2_T1         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1);
        alu3_T0         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        alu3_T1         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1);
        alu3_T2         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0);
        imm_T0          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1);
        imm_T1          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        imm_T2          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        md_T0           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0);
        md_T1           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        md_T2           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        md_T3           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1);
        branch_T0       : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1);
        branch_T1       : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        branch_T2       : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1);
        branch_T3       : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        jump_T0         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1);
        jal_T0          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        jal_T1          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1);
        in_T0           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0);
        out_T0          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        mfhi_T0         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        mflo_T0         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1);
        nop_T0          : integer := 40;
        halt_T0         : integer := 41
    );
    port(
        gra             : out    vl_logic;
        grb             : out    vl_logic;
        grc             : out    vl_logic;
        r_in            : out    vl_logic;
        r_out           : out    vl_logic;
        y_enable        : out    vl_logic;
        pc_enable       : out    vl_logic;
        mar_enable      : out    vl_logic;
        mdr_enable      : out    vl_logic;
        mdr_out         : out    vl_logic;
        ir_enable       : out    vl_logic;
        mdr_read        : out    vl_logic;
        hi_enable       : out    vl_logic;
        lo_enable       : out    vl_logic;
        zhi_enable      : out    vl_logic;
        zlo_enable      : out    vl_logic;
        inc_pc          : out    vl_logic;
        con_enable      : out    vl_logic;
        ram_enable      : out    vl_logic;
        inport_enable   : out    vl_logic;
        outport_enable  : out    vl_logic;
        inport_out      : out    vl_logic;
        pc_out          : out    vl_logic;
        zlo_out         : out    vl_logic;
        zhi_out         : out    vl_logic;
        lo_out          : out    vl_logic;
        hi_out          : out    vl_logic;
        ba_out          : out    vl_logic;
        c_out           : out    vl_logic;
        run             : out    vl_logic;
        reg_enable      : out    vl_logic_vector(15 downto 0);
        ir              : in     vl_logic_vector(31 downto 0);
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        stp             : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of r_s : constant is 1;
    attribute mti_svvh_generic_type of T0 : constant is 1;
    attribute mti_svvh_generic_type of T1 : constant is 1;
    attribute mti_svvh_generic_type of T2 : constant is 1;
    attribute mti_svvh_generic_type of T3 : constant is 1;
    attribute mti_svvh_generic_type of load_T0 : constant is 1;
    attribute mti_svvh_generic_type of load_T1 : constant is 1;
    attribute mti_svvh_generic_type of load_T2 : constant is 1;
    attribute mti_svvh_generic_type of load_T3 : constant is 1;
    attribute mti_svvh_generic_type of load_T4 : constant is 1;
    attribute mti_svvh_generic_type of loadi_T0 : constant is 1;
    attribute mti_svvh_generic_type of loadi_T1 : constant is 1;
    attribute mti_svvh_generic_type of loadi_T2 : constant is 1;
    attribute mti_svvh_generic_type of store_T0 : constant is 1;
    attribute mti_svvh_generic_type of store_T1 : constant is 1;
    attribute mti_svvh_generic_type of store_T2 : constant is 1;
    attribute mti_svvh_generic_type of store_T3 : constant is 1;
    attribute mti_svvh_generic_type of alu2_T0 : constant is 1;
    attribute mti_svvh_generic_type of alu2_T1 : constant is 1;
    attribute mti_svvh_generic_type of alu3_T0 : constant is 1;
    attribute mti_svvh_generic_type of alu3_T1 : constant is 1;
    attribute mti_svvh_generic_type of alu3_T2 : constant is 1;
    attribute mti_svvh_generic_type of imm_T0 : constant is 1;
    attribute mti_svvh_generic_type of imm_T1 : constant is 1;
    attribute mti_svvh_generic_type of imm_T2 : constant is 1;
    attribute mti_svvh_generic_type of md_T0 : constant is 1;
    attribute mti_svvh_generic_type of md_T1 : constant is 1;
    attribute mti_svvh_generic_type of md_T2 : constant is 1;
    attribute mti_svvh_generic_type of md_T3 : constant is 1;
    attribute mti_svvh_generic_type of branch_T0 : constant is 1;
    attribute mti_svvh_generic_type of branch_T1 : constant is 1;
    attribute mti_svvh_generic_type of branch_T2 : constant is 1;
    attribute mti_svvh_generic_type of branch_T3 : constant is 1;
    attribute mti_svvh_generic_type of jump_T0 : constant is 1;
    attribute mti_svvh_generic_type of jal_T0 : constant is 1;
    attribute mti_svvh_generic_type of jal_T1 : constant is 1;
    attribute mti_svvh_generic_type of in_T0 : constant is 1;
    attribute mti_svvh_generic_type of out_T0 : constant is 1;
    attribute mti_svvh_generic_type of mfhi_T0 : constant is 1;
    attribute mti_svvh_generic_type of mflo_T0 : constant is 1;
    attribute mti_svvh_generic_type of nop_T0 : constant is 1;
    attribute mti_svvh_generic_type of halt_T0 : constant is 1;
end control_unit;
