library verilog;
use verilog.vl_types.all;
entity datapath is
    port(
        pc_out          : in     vl_logic;
        zlo_out         : in     vl_logic;
        zhi_out         : in     vl_logic;
        mdr_out         : in     vl_logic;
        mdr_enable      : in     vl_logic;
        mar_enable      : in     vl_logic;
        zlo_enable      : in     vl_logic;
        zhi_enable      : in     vl_logic;
        hi_enable       : in     vl_logic;
        lo_enable       : in     vl_logic;
        hi_out          : in     vl_logic;
        lo_out          : in     vl_logic;
        c_out           : in     vl_logic;
        ram_enable      : in     vl_logic;
        pc_enable       : in     vl_logic;
        ir_enable       : in     vl_logic;
        pc_increment    : in     vl_logic;
        con_enable      : in     vl_logic;
        y_enable        : in     vl_logic;
        mdr_read        : in     vl_logic;
        gra             : in     vl_logic;
        grb             : in     vl_logic;
        grc             : in     vl_logic;
        ba_out          : in     vl_logic;
        r_in            : in     vl_logic;
        r_out           : in     vl_logic;
        outport_enable  : in     vl_logic;
        inport_enable   : in     vl_logic;
        inport_out      : in     vl_logic;
        reg_enable_in   : in     vl_logic_vector(15 downto 0);
        reg_enable_out  : in     vl_logic_vector(15 downto 0);
        opcode          : out    vl_logic_vector(4 downto 0);
        data_in         : in     vl_logic_vector(31 downto 0);
        data_inport     : in     vl_logic_vector(31 downto 0);
        data_outport    : in     vl_logic_vector(31 downto 0);
        \bus\           : out    vl_logic_vector(31 downto 0);
        clr             : in     vl_logic;
        clk             : in     vl_logic
    );
end datapath;
