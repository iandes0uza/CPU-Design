library verilog;
use verilog.vl_types.all;
entity p3_tb is
end p3_tb;
